module Sigmoid_LUT(
    input [21:0] suma,
    input predznak,
    output [15:0] vjerojatnost
);

assign vjerojatnost = (predznak!=1'b0)?(
                        (suma<22'b1001001100110011010000)?16'b0000001010001100:                             //suma veca od -4.6
                        (suma<22'b1001000000000000000000)?16'b0000001011010000:                             //suma veca od -4.5
                        (suma<22'b1000001100110011010000)?16'b0000010000101100:                             //suma veca od -4.1
                        (suma<22'b0111011001100110011000)?16'b0000011000101101:                             //suma veca od -3.7 
                        (suma<22'b0110100110011001101000)?16'b0000100100011011:                             //suma veca od -3.3 
                        (suma<22'b0101110011001100110000)?16'b0000110101011010:                             //suma veca od -2.9 
                        (suma<22'b0101000000000000000000)?16'b0001001101101011:                             //suma veca od -2.5 
                        (suma<22'b0100001100110011010000)?16'b0001101111101110:                             //suma veca od -2.1 
                        (suma<22'b0011011001100110011000)?16'b0010011110001011:                             //suma veca od -1.7 
                        (suma<22'b0010100110011001101000)?16'b0011011011010100:                             //suma veca od -1.3 
                        (suma<22'b0001110011001100110000)?16'b0100100111111111:                             //suma veca od -0.9 
                        (suma<22'b0001000000000000000000)?16'b0110000010100111:                             //suma veca od -0.5 
                        (suma<22'b0000001100110011010000)?16'b0111100110011011:16'b0000000000000000
                     ):((suma<22'b1001001100110011010000)?16'b1111110101110100:                             //suma manja od 4.6 x
                        (suma<22'b1001000000000000000000)?16'b1111110100110000:                             //suma manja od 4.5 x
                        (suma<22'b1000001100110011010000)?16'b1111101111010100:                             //suma manja od 4.1 x
                        (suma<22'b0111011001100110011000)?16'b1111100111010011:                             //suma manja od 3.7 x
                        (suma<22'b0110100110011001101000)?16'b1111011011100101:                             //suma manja od 3.3 x
                        (suma<22'b0101110011001100110000)?16'b1111001010100110:                             //suma manja od 2.9 x
                        (suma<22'b0101000000000000000000)?16'b1110110010010101:                             //suma manja od 2.5 x
                        (suma<22'b0100001100110011010000)?16'b1110010000010010:                             //suma manja od 2.1 x
                        (suma<22'b0011011001100110011000)?16'b1101100001110101:                             //suma manja od 1.7 x
                        (suma<22'b0010100110011001101000)?16'b1100100100101100:                             //suma manja od 1.3 x
                        (suma<22'b0001110011001100110000)?16'b1011011000000001:                             //suma manja od 0.9 x
                        (suma<22'b0001000000000000000000)?16'b1001111101011001:                             //suma manja od 0.5 x
                        (suma<22'b0000001100110011010000)?16'b1000011001100101:16'b1111111111111111);
endmodule